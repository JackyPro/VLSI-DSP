//=======================================
// The RCA  (4 bit)
// Design : yhchen
// Date  : 2013.3.5
// vesion : v1.0
//=======================================

module RCA4(a, b, cout, s);

    input 	[3:0]	a, b;
    output	[3:0] 	s;
    output			cout;
        
    wire	[3:0]	c;
    
    //type your design here
	//---------------------

endmodule

