`timescale 1 ns / 10 ps

module TM;

parameter 	IN_WORD_SIZE = 10;
parameter 	OUT_WORD_SIZE = 24;

reg 							clk, rst;
reg		[IN_WORD_SIZE*4-1:0] 	xin;
	

parameter   DATA_COUNT = 512*512/4;



wire	[IN_WORD_SIZE-1:0]	a0, a1, a2, a3;
wire	[OUT_WORD_SIZE-1:0]	z0, z2, z4, z6;




assign	a0 = xin[39:30];
assign	a1 = xin[29:20];
assign	a2 = xin[19:10];
assign	a3 = xin[9:0];

//===========================================//

initial
	begin
		$fsdbDumpfile("mmp.fsdb");
		$fsdbDumpvars;
	end
	
//---- gate sim -----//
//initial
//        $sdf_annotate("../mmp.sdf", U_MMP);	

//-------------------//

Top_2		U_MMP(
					.clk	(clk), 
					.rst	(rst),
					.a0		(a0),
					.a1		(a1),
					.a2		(a2),
					.a3		(a3),
					.z0		(z0),
					.z2		(z2),
					.z4		(z4),
					.z6		(z6)
				);



//*********************************
// 		control signal
//*********************************

// gen clock signal
parameter	t = 100;		
parameter	th = t/2;

always #th clk = ~clk;


initial begin
    clk = 1;
    rst = 1;
//    capture = 0;
//    mem_flag = 0;
    #th rst = 0;
    #(t*2)      rst = 1;
    #(t*10)     
	#t	xin=40'b0101000010010100010001010001110101000110;
	#t	xin=40'b0101000010010100010001010001110101000110;
	#t	xin=40'b0100111111010100011101010000010101000110;
	#t	xin=40'b0100111110010011111101001111010101000010;
	#t	xin=40'b0101000010010100001101010001000101000110;
	#t	xin=40'b0100111100010011111101001111010100111010;
	#t	xin=40'b0100111111010100001001010000100101000110;
	#t	xin=40'b0100111110010011110101010000010101000010;
	#t	xin=40'b0101000100010100010101010001010101001010;
	#t	xin=40'b0101000010010100001101010000010101000010;
	#t	xin=40'b0101000011010011111101001111010101000100;
	#t	xin=40'b0100111111010100001001010000000101000000;
	#t	xin=40'b0100110110010011011101001101100100111000;
	#t	xin=40'b0100111101010011111001001111010101000110;
	#t	xin=40'b0100111001010011110101001111000101000000;
	#t	xin=40'b0100110011010011001101001101100100110110;
	#t	xin=40'b0100111000010011011001001110100100111010;
	#t	xin=40'b0100110110010011110001001110010100111000;
	#t	xin=40'b0100111101010011101101001110100101000010;
	#t	xin=40'b0100111011010011101101001111110101000010;
	#t	xin=40'b0100110101010011100101001100100100110100;
	#t	xin=40'b0100110110010011001001001101010100111000;
	#t	xin=40'b0100110011010011011001001101000100110110;
	#t	xin=40'b0100110101010011011001001100110100111010;
	#t	xin=40'b0100110110010011011001001110000100110110;
	#t	xin=40'b0100111000010011100101001110100100111010;
	#t	xin=40'b0100110110010011010101001101100100111000;
	#t	xin=40'b0100110000010011001101001100110100110000;
	#t	xin=40'b0100110101010011010001001110000100111000;
	#t	xin=40'b0100110100010011000101001101000100110110;
	#t	xin=40'b0100110011010011001101001101010100110100;
	#t	xin=40'b0100110110010011110101001110010100111000;
	#t	xin=40'b0100110110010011100101001110000100110100;
	#t	xin=40'b0100111011010011101001001110000100111100;
	#t	xin=40'b0100110011010011011001001101000100110110;
	#t	xin=40'b0100111001010011101101001101110101000000;
	#t	xin=40'b0100111100010011110101001110110100111100;
	#t	xin=40'b0101000110010100011001010001110101001110;
	#t	xin=40'b0101000100010100010001010000100101000000;
	#t	xin=40'b0101001010010100110101010011000101001110;
	#t	xin=40'b0101001110010101000001010010110101001110;
	#t	xin=40'b0101001111010100110101010011100101001100;
	#t	xin=40'b0101001111010100111101010100000101001100;
	#t	xin=40'b0101010101010101011101010101100101011000;
	#t	xin=40'b0101011010010101011001010101110101010110;
	#t	xin=40'b0101011101010101101101010111100101100000;
	#t	xin=40'b0101011011010101101001010111100101011100;
	#t	xin=40'b0101010110010101100101010101100101010110;
	#t	xin=40'b0101010111010101100101010101100101011000;
	#t	xin=40'b0101011011010101100101010111000101011000;
	#t	xin=40'b0101010010010101000101010100110101010000;
	#t	xin=40'b0101011100010101011101010110100101011110;
	#t	xin=40'b0101001111010101000001010100010101010010;
	#t	xin=40'b0101001011010100110101010011100101001110;
	#t	xin=40'b0101000101010100000101010000000101000100;
	#t	xin=40'b0100111011010011111001010000000101000010;
	#t	xin=40'b0100101011010010100101001010110100101010;
	#t	xin=40'b0100101100010010100001001010010100101010;
	#t	xin=40'b0100100011010010011001001010110100110110;
	#t	xin=40'b0100010010010001000001000011110100011010;
	#t	xin=40'b0011111110001111110000111111010100000100;
	#t	xin=40'b0011110000001111010100111011110011101110;
	#t	xin=40'b0011101000001110000100111001010011101100;
	#t	xin=40'b0011011000001101010100110110000011010100;
	#t	xin=40'b0010111111001100001000110001110011000010;
	#t	xin=40'b0011000000001100010000110000100011000100;
	#t	xin=40'b0010111000001011011100101110100010111100;
	#t	xin=40'b0010110000001011110000101111000010111010;
	#t	xin=40'b0010101111001011001100101100100010110000;
	#t	xin=40'b0010111000001100010100110000010011000100;
	#t	xin=40'b0010111111001100001100110001110011001110;
	#t	xin=40'b0010111101001100001100110000010011000000;
	#t	xin=40'b0011000011001100100000110011000011001110;
	#t	xin=40'b0011001000001100010000110010100011001000;
	#t	xin=40'b0011001001001100100000110010100011010000;
	#t	xin=40'b0011001100001101000000110011010011010010;
	#t	xin=40'b0011010011001101001100110101100011010100;
	#t	xin=40'b0011010111001101011000110100010011010010;
	#t	xin=40'b0011010010001101011100110100100011010000;
	#t	xin=40'b0011011011001101011000110110000011011100;
	#t	xin=40'b0011011000001101010000110101110011011100;
	#t	xin=40'b0011010100001100111100110101110011011000;
	#t	xin=40'b0011010010001101010100110101110011010110;
	#t	xin=40'b0011001110001101000000110100100011010010;
	#t	xin=40'b0011001011001101001000110011000011010000;
	#t	xin=40'b0011010111001101010000110110000011011100;
	#t	xin=40'b0011010111001101011100110101010011011010;
	#t	xin=40'b0011011010001101010000110110100011011100;
	#t	xin=40'b0011010010001101000000110110000011011000;
	#t	xin=40'b0011010100001101010000110100100011011000;
	#t	xin=40'b0011010010001101001100110101010011010110;
	#t	xin=40'b0011001111001101100000110101000011011000;
	#t	xin=40'b0011011010001101101100110110010011011110;
	#t	xin=40'b0011010100001101100100110110010011011010;
	#t	xin=40'b0011010100001101000000110101000011010110;
	#t	xin=40'b0011011000001101100000110100110011011010;
	#t	xin=40'b0011010100001101010100110110100011011010;
	#t	xin=40'b0011010101001101100000110101100011011100;
	#t	xin=40'b0011011001001101100100110111010011011100;
	#t	xin=40'b0011010110001101010000110101000011011000;
	#t	xin=40'b0011010010001100111000110100010011010000;
	#t	xin=40'b0011010011001101000000110101010011010100;
	#t	xin=40'b0011010110001101110100110110010011010100;
	#t	xin=40'b0011010101001101001100110101000011011000;
	#t	xin=40'b0011011010001101100000110110100011011010;
	#t	xin=40'b0011011110001101101000110111100011011110;
	#t	xin=40'b0011100101001110001100111000110011101010;
	#t	xin=40'b0011011101001101111000110111110011011100;
	#t	xin=40'b0011100011001110101100111010010011100100;
	#t	xin=40'b0011101001001110111000111010100011101100;
	#t	xin=40'b0011101110001110110100111100000011110100;
	#t	xin=40'b0011101110001110111100111011110011101110;
	#t	xin=40'b0011101010001110010100111010000011100000;
	#t	xin=40'b0011110101001111001100111101010011110110;
	#t	xin=40'b0011110110001111000100111100000011110010;
	#t	xin=40'b0011110111001111011000111100110011110100;
	#t	xin=40'b0011111011001111110100111110010011111010;
	#t	xin=40'b0011111010001111010000111101000011110100;
	#t	xin=40'b0011111000001111010100111100110011110010;
	#t	xin=40'b0011111000001111011100111111000011111000;
	#t	xin=40'b0011111101001111101000111110100011111010;
	#t	xin=40'b0100000001010000000000111111010100000110;
	#t	xin=40'b0011111101001111101001000000000100000100;
	#t	xin=40'b0011110101001111100100111110100011110110;
	#t	xin=40'b0011111100001111011100111110000011110110;
	#t	xin=40'b0011110111001111101000111110110011111110;
	#t	xin=40'b0100000000010000011001000000100100001010;
	#t	xin=40'b0100000010010000100001000000000100000110;
	#t	xin=40'b0100000100010000100101000001110100001000;
	#t	xin=40'b0100000101010000001001000001100100000010;
	#t	xin=40'b0100000110010000100001000010100100001110;
	#t	xin=40'b0100000010010000001101000000100100000010;
	#t	xin=40'b0100000010010000011001000001100100000000;
	#t	xin=40'b0100000010010000101001000001100100000110;
	#t	xin=40'b0100000100010000000101000001010100000110;
	#t	xin=40'b0100000011010000000100111111110100000000;
	#t	xin=40'b0100001000010000010101000010110100001110;
	#t	xin=40'b0100001011010000111101000011010100010000;
	#t	xin=40'b0100000111010000010101000001010100001010;
	#t	xin=40'b0100001010010000101001000001100100001100;
	#t	xin=40'b0100000010010000100101000010110100001000;
	#t	xin=40'b0100000111010000010101000001100100000110;
	#t	xin=40'b0100000110010000000101000000110100000000;
	#t	xin=40'b0100000001001111110101000001110100000100;
	#t	xin=40'b0100001010010000101001000010100100001100;
	#t	xin=40'b0100000100001111110000111111000011111100;
	#t	xin=40'b0100000110010000011001000000010100000010;
	#t	xin=40'b0100000100010000010001000000000011111100;
	#t	xin=40'b0100001000010000100001000001110100001010;
	#t	xin=40'b0100001001010000010101000010000100000110;
	#t	xin=40'b0100000100010000010001000001000100000010;
	#t	xin=40'b0100000110010000001001000001100100000110;
	#t	xin=40'b0100000100001111111001000000000100000000;
	#t	xin=40'b0100000110010000101001000001100100001000;
	#t	xin=40'b0100000100010000010101000001000100000010;
	#t	xin=40'b0100000010010000000001000000100100000000;
	#t	xin=40'b0100001101010000100101000100000100001110;
	#t	xin=40'b0100001011010000100001000011010100001100;
	#t	xin=40'b0100001000010000101001000011110100010000;
	#t	xin=40'b0100001001010000100001000010110100001100;
	#t	xin=40'b0100000010010000011101000000100100000000;
	#t	xin=40'b0100001010010000101001000011100100001110;
	#t	xin=40'b0100000110010000110001000010010100000110;
	#t	xin=40'b0100001011010000111001000100000100001110;
	#t	xin=40'b0100001010010000110101000011000100001010;
	#t	xin=40'b0100001100010000101101000100000100001100;
	#t	xin=40'b0100001100010000111001000100000100001100;
	#t	xin=40'b0100001100010000110001000011110100001110;
	#t	xin=40'b0100001011010000100001000010100100001000;
	#t	xin=40'b0100001011010000110101000011010100001110;
	#t	xin=40'b0100000100010000100101000010000100000110;
	#t	xin=40'b0100001011010000110101000100010100010010;
	#t	xin=40'b0100001100010000110101000011010100001110;
	#t	xin=40'b0100001101010000110001000011100100001010;
	#t	xin=40'b0100001100010001000001000011100100001100;
	#t	xin=40'b0100001010010000100101000010100100001100;
	#t	xin=40'b0100001100010000111001000011110100010010;
	#t	xin=40'b0100001001010000110001000010110100001010;
	#t	xin=40'b0100001000010000100101000100000100001100;
	#t	xin=40'b0100001001010000101001000011000100001100;
	#t	xin=40'b0100001000010000101001000010000100001000;
	#t	xin=40'b0100001011010000100001000010010100001010;
	#t	xin=40'b0100001000010000100101000000110100000110;
	#t	xin=40'b0100001000010000001101000010010100001000;
	#t	xin=40'b0100000110010000101001000011010100001010;
	#t	xin=40'b0100001010010000100001000001110100001110;
	#t	xin=40'b0100001111010000101001000011010100010010;
	#t	xin=40'b0100001011010000100101000011000100001110;
	#t	xin=40'b0100001001010000100101000010010100001100;
	#t	xin=40'b0100000101010000011001000001100100000110;
	#t	xin=40'b0100001010010000101101000010110100001100;
	#t	xin=40'b0100001001010000001001000010010100000110;
	#t	xin=40'b0100001001010000111001000011010100001110;
	#t	xin=40'b0100001111010000111001000011010100010000;
	#t	xin=40'b0100000110010000110001000010100100001010;
	#t	xin=40'b0100001101010000110101000011010100001110;
	#t	xin=40'b0100001100010000110101000011010100010000;
	#t	xin=40'b0100001101010000110101000011110100010010;
	#t	xin=40'b0100001001010000101101000010010100001010;
	#t	xin=40'b0100010001010000110101000011000100010100;
	#t	xin=40'b0100001100010001000001000011100100010000;
	#t	xin=40'b0100001001010000110101000011010100001110;
	#t	xin=40'b0100001000010000101001000011100100001100;
	#t	xin=40'b0100001011010000110001000011010100010000;
	#t	xin=40'b0100000111010000110101000010110100001110;
	#t	xin=40'b0100001110010000100001000011010100010000;
	#t	xin=40'b0100001001010000101001000010000100001000;
	#t	xin=40'b0100000100010000101001000011100100001010;
	#t	xin=40'b0100010101010001010001000100000100011000;
	#t	xin=40'b0100001110010000101001000010100100001000;
	#t	xin=40'b0100000100010000011001000010100100000110;
	#t	xin=40'b0100001101010001010001000101010100010110;
	#t	xin=40'b0100010010010000101101000001100100001100;
	#t	xin=40'b0100001100010000111001000010000100001000;
	#t	xin=40'b0100000110010000010001000000100100000100;
	#t	xin=40'b0100000110010000000101000001010100001000;
	#t	xin=40'b0100001101010000100101000001010100001000;
	#t	xin=40'b0100000010010000001000111111110011111110;
	#t	xin=40'b0100000110010000010001000000110100000110;
	#t	xin=40'b0100000111010000001001000010010100001000;
	#t	xin=40'b0100001000010000100001000010000100001010;
	#t	xin=40'b0100000101010000100101000001100100000110;
	#t	xin=40'b0100000010010000000101000000110100000010;
	#t	xin=40'b0100000101010000010001000010000100001000;
	#t	xin=40'b0100000011010000011001000001110100000110;
	#t	xin=40'b0100000010010000001101000000000100000010;
	#t	xin=40'b0100001111010000110001000001010100001110;
	#t	xin=40'b0100001110010000100101000010000100001010;
	#t	xin=40'b0100000111010000110101000010010100001010;
	#t	xin=40'b0100001100010001001001000100100100010000;
	#t	xin=40'b0100000110010000010001000001000100000110;
	#t	xin=40'b0100000110010000010100111111110100001000;
	#t	xin=40'b0100000101010000011101000001100100001000;
	#t	xin=40'b0100001000010000011101000001100100001000;
	#t	xin=40'b0100000001010000010001000000110100000110;
	#t	xin=40'b0100000010010000001101000001110100001010;
	#t	xin=40'b0100000011010000010101000001010100000100;
	#t	xin=40'b0100000111010000011101000000110100000110;
	#t	xin=40'b0100001001010000100001000001010100001000;
	#t	xin=40'b0100000110010000100101000011010100001010;
	#t	xin=40'b0100001110010000110001000010100100010000;
	#t	xin=40'b0100001100010000110001000010110100001100;
	#t	xin=40'b0100001010010000011101000010000100001010;
	#t	xin=40'b0100001101010000111001000011100100001110;
	#t	xin=40'b0100001010010000100001000010000100001000;
	#t	xin=40'b0100001101010000111001000010110100001110;
	#t	xin=40'b0100001011010000101101000011010100001100;
	#t	xin=40'b0100001010010000101001000011010100010110;
	#t	xin=40'b0100000111010000100001000001110100001000;
	#t	xin=40'b0100001001010000101001000010100100001000;
	#t	xin=40'b0100001001010000100001000001100100001010;
	#t	xin=40'b0100000100010000011101000010010100001100;
	#t	xin=40'b0100000011010000010101000000110100000010;
	#t	xin=40'b0100001000010000100101000001010100000010;
	#t	xin=40'b0100001011010000100101000011000100001100;
	#t	xin=40'b0100001110010000110001000011000100010100;
	#t	xin=40'b0100010000010000111001000011110100010110;
	#t	xin=40'b0100010111010001011001000101110100011110;
	#t	xin=40'b0100001001010000110001000011000100001100;
	#t	xin=40'b0100001000010000100001000010100100001000;
	#t	xin=40'b0100000111010000101001000010000100001000;
	#t	xin=40'b0100000110010000001101000000110100000010;
	#t	xin=40'b0100000100010000001001000001010100000010;
	#t	xin=40'b0100000011010000000000111111100100000010;
	#t	xin=40'b0100000100010000011001000010010100001000;
	#t	xin=40'b0100000100010000001101000001100100001100;
	#t	xin=40'b0100000000010000001001000001010100000010;
	#t	xin=40'b0100000100010000000001000001000100000110;
	#t	xin=40'b0100000111010000010001000001010100001100;
	#t	xin=40'b0100000101010000011001000001100100001010;
	#t	xin=40'b0100001010010000011101000001010100000110;
	#t	xin=40'b0100000010010000001101000001100100000000;
	#t	xin=40'b0100000001010000000101000000100100000100;
	#t	xin=40'b0100000000001111101100111111110011111110;
	#t	xin=40'b0100000011010000011101000001110100000110;
	#t	xin=40'b0100000011010000011001000001100100001000;
	#t	xin=40'b0011111011001111111000111111100011111100;
	#t	xin=40'b0100000101010000010001000001000100000110;
	#t	xin=40'b0100001001010000010101000011010100001110;
	#t	xin=40'b0100000111010000010101000010100100001100;
	#t	xin=40'b0100000001010000001000111111110100000110;
	#t	xin=40'b0011111111001111111100111110010011111110;
	#t	xin=40'b0011111011001111110100111110100011111100;
	#t	xin=40'b0100001000010000001001000001000100000110;
	#t	xin=40'b0100000001010000000001000001010100000000;
	#t	xin=40'b0100000110010000011001000000100100000110;
	#t	xin=40'b0100001010010000110001000010100100001100;
	#t	xin=40'b0011111111001111110101000000010011111110;
	#t	xin=40'b0011111111010000001000111111010011111100;
	#t	xin=40'b0100001000010000010101000000110100001010;
	#t	xin=40'b0100000101010000010101000001100100000110;
	#t	xin=40'b0100000010010000000001000000110100000000;
	#t	xin=40'b0100000101010000001001000001010100000110;
	#t	xin=40'b0100000011010000000101000001010100000000;
	#t	xin=40'b0100000010010000001001000000110100001000;
	#t	xin=40'b0011111111001111110100111111000011111010;
	#t	xin=40'b0100000000010000000100111111010011111110;
	#t	xin=40'b0100000100010000001101000001100100000100;
	#t	xin=40'b0011111010001111111000111111000011111010;
	#t	xin=40'b0011111111001111111101000000000011111110;
	#t	xin=40'b0011111110001111111100111111100011111110;
	#t	xin=40'b0100000001001111111101000000110100001000;
	#t	xin=40'b0100000000001111101100111111000011111100;
	#t	xin=40'b0011111101001111110000111111110100000010;
	#t	xin=40'b0011111000001111011000111101100011110100;
	#t	xin=40'b0011110110001111011000111101010011111000;
	#t	xin=40'b0011110100001111100000111101100011111000;
	#t	xin=40'b0011101111001111010000111101010011110100;
	#t	xin=40'b0011101101001111001000111100110011101110;
	#t	xin=40'b0011110100001111101000111101110011110110;
	#t	xin=40'b0011110010001111000100111100010011110100;
	#t	xin=40'b0011101011001110101100111010110011101110;
	#t	xin=40'b0011101101001110101100111010010011101100;
	#t	xin=40'b0011100101001110010000111001110011100110;
	#t	xin=40'b0011100001001101111100111001100011100000;
	#t	xin=40'b0011100101001110000000110111100011100010;
	#t	xin=40'b0011100010001110000100111000100011100110;
	#t	xin=40'b0011010100001101000000110100100011010010;
	#t	xin=40'b0011010001001100111000110100010011001110;
	#t	xin=40'b0011010100001100111100110011110011001110;
	#t	xin=40'b0011001011001100111000110011010011010000;
	#t	xin=40'b0011010101001101011000110111100011100000;
	#t	xin=40'b0011100111001110011100111000100011101010;
	#t	xin=40'b0011101010001110110100111011100011101100;
	#t	xin=40'b0011110100001111010000111101000011110100;
	#t	xin=40'b0011111111010000001001000001000100001000;
	#t	xin=40'b0100000110010000010001000001110100001110;
	#t	xin=40'b0100010101010001000001000101110100011000;
	#t	xin=40'b0100010110010001010001000101010100011000;
	#t	xin=40'b0100011101010001110001001000000100100000;
	#t	xin=40'b0100100001010010001101001000110100100100;
	#t	xin=40'b0100100111010010110001001011010100101100;
	#t	xin=40'b0100101101010010101001001100000100110010;
	#t	xin=40'b0100110100010010111001001011010100110000;
	#t	xin=40'b0100110010010011010001001100110100110100;
	#t	xin=40'b0100111001010011110101001110110100111110;
	#t	xin=40'b0100111010010011110101001111000100111110;
	#t	xin=40'b0100111100010011110101010000000100111110;
	#t	xin=40'b0101000001010100000101010000100101000110;
	#t	xin=40'b0101000001010011110101010000100100111100;
	#t	xin=40'b0101000100010100011001010000100101000110;
	#t	xin=40'b0101000001010011111101001111110101000010;
	#t	xin=40'b0100111011010011011001001110100100110110;
	#t	xin=40'b0100110111010011011101001101010100111000;
	#t	xin=40'b0100110011010010111101001011010100101000;
	#t	xin=40'b0100110010010010111001001011100100101100;
	#t	xin=40'b0100110000010011001101001100110100110100;
	#t	xin=40'b0100101110010010111101001100000100101100;
	#t	xin=40'b0100110000010011001001001100100100110100;
	#t	xin=40'b0100101110010011000001001011100100101110;
	#t	xin=40'b0100110010010011000001001100100100101110;
	#t	xin=40'b0100110100010011001101001100100100110110;
	#t	xin=40'b0100101011010010111101001010010100101110;
	#t	xin=40'b0100110110010011010001001101100100111010;
	#t	xin=40'b0100110101010011100101001101110100110110;
	#t	xin=40'b0100110001010011000101001011000100110000;
	#t	xin=40'b0100110111010011101101001101110100111010;
	#t	xin=40'b0100110100010011001001001110000100111000;
	#t	xin=40'b0100110100010011010001001100100100110100;
	#t	xin=40'b0100110001010011001001001100110100110100;
	#t	xin=40'b0100111011010011111001001110010101000000;
	#t	xin=40'b0100110110010011100101001101010100111100;
	#t	xin=40'b0100110100010011011001001101110100110110;
	#t	xin=40'b0100111110010011100001001110100100111010;
	#t	xin=40'b0100110110010011010001001101010100110100;
	#t	xin=40'b0100110011010011001101001101000100110100;
	#t	xin=40'b0100110011010011000101001100010100101110;
	#t	xin=40'b0100111000010011010101001101100100111100;
	#t	xin=40'b0100110101010011001101001100100100110010;
	#t	xin=40'b0100110001010011000001001100010100101110;
	#t	xin=40'b0100110011010011001001001100010100110100;
	#t	xin=40'b0100110011010011001001001100000100110010;
	#t	xin=40'b0100110100010011001001001101000100110110;
	#t	xin=40'b0100101111010011010001001100010100110010;
	#t	xin=40'b0100110001010011010001001100010100110000;
	#t	xin=40'b0100110010010011011001001101010100110010;
	#t	xin=40'b0100110100010011010101001100000100110010;
	#t	xin=40'b0100110010010011001101001100100100101110;
	#t	xin=40'b0100110000010011001101001011110100110000;
	#t	xin=40'b0100111001010011011101001110010100111100;
	#t	xin=40'b0100110110010011010001001110000100110100;
	#t	xin=40'b0100110001010011001101001110010100110100;
	#t	xin=40'b0100110000010011000101001101000100110010;
	#t	xin=40'b0100101111010011000001001100010100110000;
	#t	xin=40'b0100110011010011010001001101000100110100;
	#t	xin=40'b0100110101010011011001001110100100111100;
	#t	xin=40'b0100110101010011010001001100100100110100;
	#t	xin=40'b0100110110010011110101001110010100111110;
	#t	xin=40'b0100111001010011100101001110100100111100;
	#t	xin=40'b0100110111010011011101001110110100111010;
	#t	xin=40'b0100110010010011011101001101010100110100;
	#t	xin=40'b0100110101010011011001001101110100110110;
	#t	xin=40'b0100111100010011100001001110110100111000;
	#t	xin=40'b0100111101010011100001001110010101000000;
	#t	xin=40'b0100111100010011101101001110100100111110;
	#t	xin=40'b0100111100010011110001001111000100111110;
	#t	xin=40'b0100111001010011011101001110100100111010;
	#t	xin=40'b0100110110010011100001001110000100111000;
	#t	xin=40'b0100111001010011011101001101100100111000;
	#t	xin=40'b0100110001010011001001001100010100110000;
	#t	xin=40'b0100110111010011010001001100100100111000;
	#t	xin=40'b0100110011010011000101001100110100110110;
	#t	xin=40'b0100110011010011011001001110110100111100;
	#t	xin=40'b0101000111010101001101010110110101100010;
	#t	xin=40'b0101100110010111000001011110110110000010;
	#t	xin=40'b0101111100011000100001100010010110001110;
	#t	xin=40'b0110010000011001010101100101100110011100;
	#t	xin=40'b0110011010011001110001101000000110100000;
	#t	xin=40'b0110100010011010011001101010000110101010;
	#t	xin=40'b0110100101011010101001101010100110101010;
	#t	xin=40'b0110101001011010101001101011000110101010;
	#t	xin=40'b0110101111011010111101101011110110110000;
	#t	xin=40'b0110110001011011001101101100100110110100;
	#t	xin=40'b0110110011011011010001101101100110110110;
	#t	xin=40'b0110110011011011010001101101000110110100;
	#t	xin=40'b0110110100011011011001101101000110110100;
	#t	xin=40'b0110110110011011100001101101100110111000;
	#t	xin=40'b0110110010011011001101101101000110110000;
	#t	xin=40'b0110101101011010110001101010110110100110;
	#t	xin=40'b0110100011011010000001100111010110011000;
	#t	xin=40'b0110010010011000111001100010000110000000;
	#t	xin=40'b0101110101010111000001011001110101011000;
	#t	xin=40'b0101010011010100101101001111000100110000;
	#t	xin=40'b0100100011010001010101000001100011110100;
	#t	xin=40'b0011110110001110101100110110010011010100;
	#t	xin=40'b0011100100001101010100110011110011010010;
	#t	xin=40'b0011001011001100111000110001100011001010;
	#t	xin=40'b0011001000001100101000110011110011001110;
	#t	xin=40'b0011001111001100111000110011100011010000;
	#t	xin=40'b0011010111001101011000110110000011011110;
	#t	xin=40'b0011011001001101011000110110100011010010;
	#t	xin=40'b0011011101001101101000111000000011100010;
	#t	xin=40'b0011100110001110010100111000110011101000;
	#t	xin=40'b0011100111001110101000111011100011101010;
	#t	xin=40'b0011101101001110110000111011000011110000;
	#t	xin=40'b0011101001001110100100111011010011101100;
	#t	xin=40'b0011101101001110111100111011000011101110;
	#t	xin=40'b0011101110001111001000111011000011101100;
	#t	xin=40'b0011101011001110111100111100010011110010;
	#t	xin=40'b0011110000001110111100111101100011111000;
	#t	xin=40'b0011110111001111011100111110000011111110;
	#t	xin=40'b0011101110001111010000111101110011110010;
	#t	xin=40'b0011101110001111000000111100010011101110;
	#t	xin=40'b0011101110001110110000111100000011101100;
	#t	xin=40'b0011110001001111000100111011010011110000;
	#t	xin=40'b0011110001001111011100111110000011111010;
	#t	xin=40'b0011110101001111100000111100110011110010;
	#t	xin=40'b0011101101001111000000111100100011101100;
	#t	xin=40'b0011110001001111010100111101100011110110;
	#t	xin=40'b0011110011001111011000111101100011110100;
	#t	xin=40'b0011111001001111101000111110000011111010;
	#t	xin=40'b0011111011001111111000111110100100000000;
	#t	xin=40'b0011110111001111000100111100100011110010;
	#t	xin=40'b0011110001001111000000111101000011110000;
	#t	xin=40'b0011111010001111001000111100100011111000;
	#t	xin=40'b0011110011001110111100111011010011101100;
	#t	xin=40'b0011110100001111010100111011100011110010;
	#t	xin=40'b0011111000001111010000111101110011110110;
	#t	xin=40'b0011110011001111100000111101000011111000;
	#t	xin=40'b0011110010001111000000111011000011101110;
	#t	xin=40'b0011110101001111100100111101010011110110;
	#t	xin=40'b0011110101001110111100111100010011110010;
	#t	xin=40'b0011111000001111001100111101000011110010;
	#t	xin=40'b0011110111001111110000111110100011110110;
	#t	xin=40'b0011110110001111011100111110000011110100;
	#t	xin=40'b0011111001001111100000111101110011111000;
	#t	xin=40'b0100000000001111110100111111100100000010;
	#t	xin=40'b0011110100001111011000111101000011101110;
	#t	xin=40'b0011110110001111101100111110110011111000;
	#t	xin=40'b0011111110001111011000111110000011111100;
	#t	xin=40'b0011111010001111101000111101010011111010;
	#t	xin=40'b0011110111001111100100111111000011111100;
	#t	xin=40'b0011111011001111101000111111100011111100;
	#t	xin=40'b0011111010001111100100111110110011111110;
	#t	xin=40'b0011110010001111001000111101100011110110;
	#t	xin=40'b0011111010001111110000111111010011111000;
	#t	xin=40'b0011111000001111101000111110010011111010;
	#t	xin=40'b0011110110001111100000111110000011111010;
	#t	xin=40'b0011110100001111001100111011000011101100;
	#t	xin=40'b0011101111001111000000111011000011101100;
	#t	xin=40'b0011111011001111110001000000000100000010;
	#t	xin=40'b0011110001001111010100111101000011110100;
	#t	xin=40'b0011111010001111111000111110000011111110;
	#t	xin=40'b0011111101001111100100111110110011111100;
	#t	xin=40'b0011111101001111101100111111110011111100;
	#t	xin=40'b0100000010010000000101000000010100000100;
	#t	xin=40'b0011111110001111010100111110110011111000;
	#t	xin=40'b0011111111001111100100111110110011111110;
	#t	xin=40'b0011110110001111100000111111000011111010;
	#t	xin=40'b0011111000001111011000111101110011110010;
	#t	xin=40'b0100000010001111111001000000100100000010;
	#t	xin=40'b0011111111001111110000111110100011111010;
	#t	xin=40'b0011111110001111101100111110100011111100;
	#t	xin=40'b0011111111001111110100111111000011111110;
	#t	xin=40'b0011110101001111011100111100010011110000;
	#t	xin=40'b0011111001001111011100111101110011110110;
	#t	xin=40'b0011101101001110101000111010010011100100;
	#t	xin=40'b0011110110001111001000111011000011110010;
	#t	xin=40'b0011101100001110101000111001100011101000;
	#t	xin=40'b0011110111001111011000111100100011101110;
	#t	xin=40'b0011110111001111010000111100000011101100;
	#t	xin=40'b0011110001001111000100111011010011100110;
	#t	xin=40'b0011111000001111101100111101110011110010;
	#t	xin=40'b0011111000001111111000111110110011111000;
	#t	xin=40'b0011111100010000100101000101000100010100;
	#t	xin=40'b0100000011010010010001001100110101001000;
	#t	xin=40'b0011111011010010001001001111100101010000;
	#t	xin=40'b0011110000010001101001001111000101010100;
	#t	xin=40'b0011101111010000100101001101110101011000;
	#t	xin=40'b0011011100001111100101001001100101010100;
	#t	xin=40'b0011010010001101101101000000100100110110;
	#t	xin=40'b0010101111001011101100110011010100000000;
	#t	xin=40'b0100111001010011100101001110010100111010;
	#t	xin=40'b0100111001010011100101001110010100111010;
	#t	xin=40'b0100111110010011110101001110100100111010;
	#t	xin=40'b0100111011010011101001001111100100111011;
	#t	xin=40'b0100111011010011011001001111100100111100;
	#t	xin=40'b0100111110010011100101001110000100110101;
	#t	xin=40'b0100111010010011100101001101110100110110;
	#t	xin=40'b0100111000010011101001001101000100110001;
	#t	xin=40'b0101000001010011110101001111010100111111;
	#t	xin=40'b0100111011010011011101001110100100111010;
	#t	xin=40'b0100111011010011010001001110000100111100;
	#t	xin=40'b0100111111010011110001001110100100111001;
	#t	xin=40'b0100111011010011101101001110110100111000;
	#t	xin=40'b0100110110010011101001001101010100110100;
	#t	xin=40'b0100110110010011100101001110000100111010;
	#t	xin=40'b0100111001010011001101001110110100111011;
	#t	xin=40'b0100111001010011011101001111000100111000;
	#t	xin=40'b0100110110010011101001001110010100111100;
	#t	xin=40'b0100111111010011010001001101110101000001;
	#t	xin=40'b0100111100010011010101001101100100110011;
	#t	xin=40'b0100111001010011010001001111010100111010;
	#t	xin=40'b0100110101010011100101001111000100111001;
	#t	xin=40'b0100110110010011011001001100110100111010;
	#t	xin=40'b0100110100010011001101001101100100111000;
	#t	xin=40'b0100110100010011001001001100110100110011;
	#t	xin=40'b0100110110010011100001001101000100110010;
	#t	xin=40'b0100101111010011001001001100100100110010;
	#t	xin=40'b0100111001010011011001001101110100110110;
	#t	xin=40'b0100101111010011010101001101100100110110;
	#t	xin=40'b0100110100010011000101001111000100110110;
	#t	xin=40'b0100111011010011011101001101000100110001;
	#t	xin=40'b0100111011010011101101001101000100110110;
	#t	xin=40'b0100111111010011100101001110000100110101;
	#t	xin=40'b0100111100010011011001001110110100111001;
	#t	xin=40'b0100111100010100000001001110110101000001;
	#t	xin=40'b0101000011010100100101010001000101000010;
	#t	xin=40'b0101001010010100101101010001100101001001;
	#t	xin=40'b0101000101010100100101010001110101000101;
	#t	xin=40'b0101010001010100111001010011100101001011;
	#t	xin=40'b0101001110010100110101010011100101010010;
	#t	xin=40'b0101010101010101001001010101010101010001;
	#t	xin=40'b0101010011010101000001010011100101010001;
	#t	xin=40'b0101011100010101001001010011100101010100;
	#t	xin=40'b0101010000010101000101010101010101010100;
	#t	xin=40'b0101010010010101001001010110000101010101;
	#t	xin=40'b0101010010010101100001010101110101010000;
	#t	xin=40'b0101010001010101001001010101010101010010;
	#t	xin=40'b0101011000010101001101010100000101011010;
	#t	xin=40'b0101010110010101010101010100000101010011;
	#t	xin=40'b0101001001010101001001010100110101010110;
	#t	xin=40'b0101001101010100111001010010110101010001;
	#t	xin=40'b0101001010010100111101010010110101001101;
	#t	xin=40'b0101000101010100110101010001110101001110;
	#t	xin=40'b0101000000010011110001010000100101001010;
	#t	xin=40'b0100111011010011100101001111000100111111;
	#t	xin=40'b0100101111010011001001001010010100101001;
	#t	xin=40'b0100100010010010011101001001000100011111;
	#t	xin=40'b0100100011010001111001000110110100010111;
	#t	xin=40'b0100001110010001001101000011110100010001;
	#t	xin=40'b0100001010010000011101000100010100000111;
	#t	xin=40'b0011110101001111011100111111110011111100;
	#t	xin=40'b0011101100001111100000111011110011101001;
	#t	xin=40'b0011011101001110001000110111110011010111;
	#t	xin=40'b0011100011001101010100110100010011010001;
	#t	xin=40'b0011000110001100010100110010000011000100;
	#t	xin=40'b0010111011001011101000101101010010111011;
	#t	xin=40'b0010110111001011100100101100010010101101;
	#t	xin=40'b0010110000001011010100101101000010110101;
	#t	xin=40'b0010110100001011001000101110110010101111;
	#t	xin=40'b0010111001001011101100101101110010101111;
	#t	xin=40'b0010111000001011101000101110110010111000;
	#t	xin=40'b0010111010001011100000101111000010111101;
	#t	xin=40'b0010111010001100000000110001110010111011;
	#t	xin=40'b0011001000001100000000110000100010111101;
	#t	xin=40'b0011001011001100100100110001100011000011;
	#t	xin=40'b0011001111001100111000110010100011001010;
	#t	xin=40'b0011010010001100100000110010100011000101;
	#t	xin=40'b0011001100001100010000110001110011001011;
	#t	xin=40'b0011010000001100110100110101000011010011;
	#t	xin=40'b0011001101001100111100110100010011001111;
	#t	xin=40'b0011010100001101001100110100010011001101;
	#t	xin=40'b0011011001001101000100110011100011001101;
	#t	xin=40'b0011011010001101010100110101100011010010;
	#t	xin=40'b0011001111001101001100110101110011010011;
	#t	xin=40'b0011010100001100101000110100100011010000;
	#t	xin=40'b0011010000001101010100110100110011010111;
	#t	xin=40'b0011010110001101011100110100010011010111;
	#t	xin=40'b0011010101001101101000110100100011010111;
	#t	xin=40'b0011001011001101001000110101110011010111;
	#t	xin=40'b0011010010001101101100110110000011010000;
	#t	xin=40'b0011010101001101010100110101100011010011;
	#t	xin=40'b0011010001001101001100110100110011001101;
	#t	xin=40'b0011010100001100111100110011000011001101;
	#t	xin=40'b0011010000001100101100110011100011001000;
	#t	xin=40'b0011010110001101000000110100100011010100;
	#t	xin=40'b0011001111001101000000110011100011001111;
	#t	xin=40'b0011010010001101000000110011010011001101;
	#t	xin=40'b0011011000001101000100110011010011010101;
	#t	xin=40'b0011011001001100110100110011010011010001;
	#t	xin=40'b0011001011001100011000110011000011001011;
	#t	xin=40'b0011001111001100101000110101000011001011;
	#t	xin=40'b0011010011001101001000110101000011001100;
	#t	xin=40'b0011010010001101001100110101010011010001;
	#t	xin=40'b0011011111001101011100110111100011010111;
	#t	xin=40'b0011011101001101110100111000010011100011;
	#t	xin=40'b0011011111001101011100110111000011011111;
	#t	xin=40'b0011011100001101100100110111000011011110;
	#t	xin=40'b0011011111001110010000110111100011100101;
	#t	xin=40'b0011011101001110010000111001010011100001;
	#t	xin=40'b0011100011001110011100111001110011100101;
	#t	xin=40'b0011101110001110011100111011110011100110;
	#t	xin=40'b0011100110001110101000111011010011101011;
	#t	xin=40'b0011101011001110101100111100100011101011;
	#t	xin=40'b0011101110001110101100111100000011101111;
	#t	xin=40'b0011110001001111010000111100010011101101;
	#t	xin=40'b0011110100001111000000111101010011110010;
	#t	xin=40'b0011110000001111001000111101010011111010;
	#t	xin=40'b0011110101001111100000111101110011110100;
	#t	xin=40'b0011111101001111100100111100000011111010;
	#t	xin=40'b0011111000001111010100111100110011110111;
	#t	xin=40'b0011111101001111101000111101000011110101;
	#t	xin=40'b0011111100001111111000111101100011111110;
	#t	xin=40'b0100000011001111100000111101100011110110;
	#t	xin=40'b0011111010001111010100111111010100000010;
	#t	xin=40'b0011111100001111011100111110010100000001;
	#t	xin=40'b0011111101001111100000111110010011110111;
	#t	xin=40'b0100000111010000001001000000100100000000;
	#t	xin=40'b0011111111001111110100111111100011111100;
	#t	xin=40'b0011111001001111110100111110110011111011;
	#t	xin=40'b0011111101010000000001000000100100000001;
	#t	xin=40'b0011111111001111111000111111110100000010;
	#t	xin=40'b0100000000010000001000111111110011111010;
	#t	xin=40'b0100000011001111111000111110110100000010;
	#t	xin=40'b0100000001001111111001000000010011111100;
	#t	xin=40'b0100001001010000001101000000100100001110;
	#t	xin=40'b0100000011001111110101000000000011111111;
	#t	xin=40'b0100000010010000000101000001100011111110;
	#t	xin=40'b0100000100001111111001000000000100000001;
	#t	xin=40'b0100001000010000010101000001100100000100;
	#t	xin=40'b0100000001010000000001000001010100000001;
	#t	xin=40'b0100000011010000011001000001000011111111;
	#t	xin=40'b0100000111010000001001000001000100000110;
	#t	xin=40'b0011111111010000111101000010010100001110;
	#t	xin=40'b0100000111010000001001000000100100001000;
	#t	xin=40'b0100000110010000011101000001100100000111;
	#t	xin=40'b0100000011010000010001000001100100001110;
	#t	xin=40'b0100001000010000001001000010100100001000;
	#t	xin=40'b0100000101010000010001000010010100000100;
	#t	xin=40'b0100000011010000011101000011000100000100;
	#t	xin=40'b0100000111010000000101000001010100000101;
	#t	xin=40'b0100000101010000001001000000100100000011;
	#t	xin=40'b0100000100010000010001000001010100000101;
	#t	xin=40'b0100000010010000011001000000010100000100;
	#t	xin=40'b0100000011010000100001000001110100001001;
	#t	xin=40'b0100000101010000001101000000110100000100;
	#t	xin=40'b0100000000001111111101000000100100000000;
	#t	xin=40'b0100000100010000100101000001010100000000;
	#t	xin=40'b0100001100010000001001000010010100000110;
	#t	xin=40'b0100000111010000011001000011010100001100;
	#t	xin=40'b0100001100010000100101000001000100000011;
	#t	xin=40'b0100000011010000001100111111000100000000;
	#t	xin=40'b0100001100010000011101000010100100000010;
	#t	xin=40'b0100001011010000010101000010010100001100;
	#t	xin=40'b0100000110010000010101000001010100000100;
	#t	xin=40'b0100000111010000100101000010110100001100;
	#t	xin=40'b0100001100010000010101000011000100001110;
	#t	xin=40'b0100001001010000100001000010100100000110;
	#t	xin=40'b0100001011010000101001000001110100001011;
	#t	xin=40'b0100000110010000101101000001100100001000;
	#t	xin=40'b0100001000010000011101000010010100001001;
	#t	xin=40'b0100010000010000110001000010100100000101;
	#t	xin=40'b0100001110010001000101000010000100001001;
	#t	xin=40'b0100000110010001000001000011100100001001;
	#t	xin=40'b0100001010010000111001000011100100001011;
	#t	xin=40'b0100001011010000101101000010010100001101;
	#t	xin=40'b0100000101010000100101000011100100001001;
	#t	xin=40'b0100001001010000011101000001110100001001;
	#t	xin=40'b0100001000010000001001000100000100001001;
	#t	xin=40'b0100001010010000100101000011000100001011;
	#t	xin=40'b0100001000010000101001000001110100000011;
	#t	xin=40'b0100001010010001001001000000000100001000;
	#t	xin=40'b0100000110010000011001000001010100001010;
	#t	xin=40'b0100001010010000101101000000100100000101;
	#t	xin=40'b0100001001010000100101000010000100001001;
	#t	xin=40'b0100000111010000101001000010010100001011;
	#t	xin=40'b0100000010010000100001000000110100001010;
	#t	xin=40'b0100010001010000101101000010000100001000;
	#t	xin=40'b0100001110010001000101000010100100001101;
	#t	xin=40'b0100001001010000110101000010110100000001;
	#t	xin=40'b0100000100010000111001000011000100000111;
	#t	xin=40'b0100000101010000010101000010100100000111;
	#t	xin=40'b0100001001010000010101000001010100001011;
	#t	xin=40'b0100000100010000111001000000010100000110;
	#t	xin=40'b0100000111010000010101000010110100001011;
	#t	xin=40'b0100001010010000011101000001000100001001;
	#t	xin=40'b0100001101010000011101000010000100000100;
	#t	xin=40'b0100000110010000100101000001010100000111;
	#t	xin=40'b0100000110010000000101000000000100000100;
	#t	xin=40'b0100001110010000110001000010110100001001;
	#t	xin=40'b0100001100010000101101000010110100000111;
	#t	xin=40'b0100001000010000011001000010010100001011;
	#t	xin=40'b0100000101010000011000111111010100000000;
	#t	xin=40'b0100000101010000100101000010000100000110;
	#t	xin=40'b0100001001010000111001000010010100000110;
	#t	xin=40'b0100000110010000010001000010100100001010;
	#t	xin=40'b0100001001010000010101000000010100000110;
	#t	xin=40'b0100000100010000011001000010010100000100;
	#t	xin=40'b0100000110001111110101000001010100001010;
	#t	xin=40'b0100000111010000100001000001010100000110;
	#t	xin=40'b0100000000010000001101000001100100001010;
	#t	xin=40'b0100000110010000100101000010110100001111;
	#t	xin=40'b0100001010010000101001000001010100001000;
	#t	xin=40'b0100001001010000100101000011000100001000;
	#t	xin=40'b0100001010001111110001000000000100001001;
	#t	xin=40'b0100001001010000100001000001110100000100;
	#t	xin=40'b0100001011010000010101000001010100001001;
	#t	xin=40'b0100001000010000100001000001010100000101;
	#t	xin=40'b0100000011001111111100111111100100000100;
	#t	xin=40'b0100000000010000010101000001110100000101;
	#t	xin=40'b0100000100010000000101000001000100000001;
	#t	xin=40'b0011111111010000010101000000000100000100;
	#t	xin=40'b0100000001010000001001000000110100000110;
	#t	xin=40'b0100001001010000010000111111110100000100;
	#t	xin=40'b0100000010001111111000111111000100001001;
	#t	xin=40'b0100000100010000010101000001010100000001;
	#t	xin=40'b0100001011010000100000111111100100000101;
	#t	xin=40'b0100000111010000110001000000110100000110;
	#t	xin=40'b0100001001010000011101000001110100000011;
	#t	xin=40'b0100010000010000000101000001100100001001;
	#t	xin=40'b0100001000010000000001000000110100000100;
	#t	xin=40'b0100001001010000011101000000110100001010;
	#t	xin=40'b0100001001010000010101000001110100000111;
	#t	xin=40'b0100000001010000000101000001100011111111;
	#t	xin=40'b0011111110001111101100111111000100000010;
	#t	xin=40'b0100000101001111101001000000000100000001;
	#t	xin=40'b0100001000010000001101000000110100000100;
	#t	xin=40'b0100000111010000001101000001110100000010;
	#t	xin=40'b0100000111010000010001000010100100001000;
	#t	xin=40'b0100001000010000010101000000000100000100;
	#t	xin=40'b0100000101010000010001000001100100001001;
	#t	xin=40'b0100001000010000100001000100000100000101;
	#t	xin=40'b0100001001010000001001000010000100001101;
	#t	xin=40'b0100001000010000011001000010000100001100;
	#t	xin=40'b0100001100010000110101000001110100001111;
	#t	xin=40'b0100000101010000100001000100000100001011;
	#t	xin=40'b0100001010010000100001000010010100010010;
	#t	xin=40'b0100001101010000110101000001010100001010;
	#t	xin=40'b0100001100010000010001000001010100001100;
	#t	xin=40'b0100000111010000101101000011000100000101;
	#t	xin=40'b0100000011010000001001000000110100001011;
	#t	xin=40'b0100000101010000001001000000110100000100;
	#t	xin=40'b0100000011010000011101000001010100000101;
	#t	xin=40'b0100001110010000010001000010000100010001;
	#t	xin=40'b0100001110010000010101000000100011111011;
	#t	xin=40'b0100000101010000011001000000110100000100;
	#t	xin=40'b0100000011010000011101000001000100000100;
	#t	xin=40'b0100000110010000001101000001010011111111;
	#t	xin=40'b0100000100010000010101000001110100000000;
	#t	xin=40'b0100001001010001000001000001110100001010;
	#t	xin=40'b0100001000010000001101000000110100000010;
	#t	xin=40'b0100000110010000001101000001010100000110;
	#t	xin=40'b0100001010010000100101000000110100000100;
	#t	xin=40'b0100000000010000100001000010000100001101;
	#t	xin=40'b0100000011010000001001000000000100000011;
	#t	xin=40'b0100000101010000001101000001000100001000;
	#t	xin=40'b0100000010010000010101000011000100000111;
	#t	xin=40'b0100000000001111110101000000010100001001;
	#t	xin=40'b0100001001010000011001000010100100000011;
	#t	xin=40'b0100001000010000100001000001100100000001;
	#t	xin=40'b0011111101001111111000111111110100000100;
	#t	xin=40'b0100000010010000001000111111100100000100;
	#t	xin=40'b0100000101010000001101000000110100000000;
	#t	xin=40'b0011111101010000001100111111110100000011;
	#t	xin=40'b0011111111001111111000111111000100000001;
	#t	xin=40'b0100000100010000011101000010000100000000;
	#t	xin=40'b0011111010001111111000111111100100000110;
	#t	xin=40'b0011111101010000001001000000110100000100;
	#t	xin=40'b0011111111010000000000111111100100000110;
	#t	xin=40'b0100000010001111110001000000100100000010;
	#t	xin=40'b0011111110010000000001000000000100000010;
	#t	xin=40'b0011111101001111110100111111000100000000;
	#t	xin=40'b0011111111001111110101000000100011111111;
	#t	xin=40'b0011111101010000000101000000110100000100;
	#t	xin=40'b0011111101001111110000111110110100000100;
	#t	xin=40'b0100000100001111101100111111110011111110;
	#t	xin=40'b0100000011010000000001000001000011111101;
	#t	xin=40'b0100000011001111100100111111100100001100;
	#t	xin=40'b0100000100001111110101000000000011111110;
	#t	xin=40'b0011111101010000000100111111110100000000;
	#t	xin=40'b0100000011001111111100111110010011111001;
	#t	xin=40'b0100000111001111111001000000000011111110;
	#t	xin=40'b0011111110010000010000111111110011111110;
	#t	xin=40'b0100000000010000001001000001000100000001;
	#t	xin=40'b0100000001001111111001000001000100000001;
	#t	xin=40'b0100000011010000000101000000100100000010;
	#t	xin=40'b0100000011001111110100111111110100000000;
	#t	xin=40'b0100000000010000010001000000010011111100;
	#t	xin=40'b0100000000010000001101000001000011111101;
	#t	xin=40'b0100000000001111011100111111110100000011;
	#t	xin=40'b0100000101001111111101000000010011111110;
	#t	xin=40'b0011111110001111101101000001000100000010;
	#t	xin=40'b0011111110010000100001000001010100000101;
	#t	xin=40'b0100000001001111101000111111000011111111;
	#t	xin=40'b0011111011001111100100111111110011111010;
	#t	xin=40'b0011111111001111010000111111000011111010;
	#t	xin=40'b0100000010001111100100111100000011111110;
	#t	xin=40'b0011110101001111011100111101000011111010;
	#t	xin=40'b0011111110001111111100111110010011110010;
	#t	xin=40'b0011110101001111000100111010100011110001;
	#t	xin=40'b0011110000001111001000111101010011110000;
	#t	xin=40'b0011110100001111001000111100100011110100;
	#t	xin=40'b0011101100001110111100111011110011110010;
	#t	xin=40'b0011100110001110101000111010010011101001;
	#t	xin=40'b0011101000001110100100111010010011100110;
	#t	xin=40'b0011100111001110011100111000110011100011;
	#t	xin=40'b0011011011001101101100111000000011101000;
	#t	xin=40'b0011100010001110001000110111110011011110;
	#t	xin=40'b0011100101001110000100110110000011011111;
	#t	xin=40'b0011101101001101011000110111110011011100;
	#t	xin=40'b0011010101001110001100110111000011011110;
	#t	xin=40'b0011010101001101001000110111100011010011;
	#t	xin=40'b0011010111001101010000110110100011011100;
	#t	xin=40'b0011010011001101001000110100110011010011;
	#t	xin=40'b0011010011001101011100110010110011010100;
	#t	xin=40'b0011011100001101011100110100010011001111;
	#t	xin=40'b0011011111001101110100110110100011010011;
	#t	xin=40'b0011100011001110001100111000110011100000;
	#t	xin=40'b0011110100001110110100111100100011110000;
	#t	xin=40'b0011110111001111100000111110110011111000;
	#t	xin=40'b0100000000001111111001000010110100000101;
	#t	xin=40'b0100001011010000101001000011110100001010;
	#t	xin=40'b0100011011010001010101000101110100011000;
	#t	xin=40'b0100011000010001110101000111100100010110;
	#t	xin=40'b0100101010010010100001001001010100100100;
	#t	xin=40'b0100100111010010100101001001010100101001;
	#t	xin=40'b0100101100010010100101001010110100101011;
	#t	xin=40'b0100110001010011001001001101000100101110;
	#t	xin=40'b0100110101010011000101001101000100110001;
	#t	xin=40'b0100110101010011100101001110000100110010;
	#t	xin=40'b0100111001010011100001001111000100111100;
	#t	xin=40'b0101000001010011111101001111110101000011;
	#t	xin=40'b0100111100010100001101010000100100111110;
	#t	xin=40'b0100111110010100000001010001000101000001;
	#t	xin=40'b0100111011010100001001001111000100111101;
	#t	xin=40'b0100111101010100000101001111110100111101;
	#t	xin=40'b0100111100010011011101010000000100111101;
	#t	xin=40'b0100111100010100000101001110110100111101;
	#t	xin=40'b0100111101010011110001001100110100110100;
	#t	xin=40'b0100111000010011101101001110100100110100;
	#t	xin=40'b0100111011010011110001001110000100111111;
	#t	xin=40'b0100111010010011100101001101100100110111;
	#t	xin=40'b0100111001010011011101001101010100111100;
	#t	xin=40'b0100111000010011101001001110000100110011;
	#t	xin=40'b0100111001010100000101001110100100110111;
	#t	xin=40'b0100111110010011110101001110010100111010;
	#t	xin=40'b0100111101010100000001010001000100111101;
	#t	xin=40'b0100111100010011110001010000000100111101;
	#t	xin=40'b0100111101010011110001001111100100111011;
	#t	xin=40'b0100111001010100001101010000000100111010;
	#t	xin=40'b0100111011010011111101001111100100111110;
	#t	xin=40'b0100111101010100001101010000010101000000;
	#t	xin=40'b0101000000010011110001001111000101000001;
	#t	xin=40'b0100111110010011110101001111010100111100;
	#t	xin=40'b0101000000010011110101001111110100111010;
	#t	xin=40'b0100111100010011111001001110110101000000;
	#t	xin=40'b0100111011010011101101001111010100111100;
	#t	xin=40'b0100111110010011100001001111010100111001;
	#t	xin=40'b0100111101010011101001001110100100111101;
	#t	xin=40'b0100111000010011100001001101100100111011;
	#t	xin=40'b0100111101010011100101001111000100111101;
	#t	xin=40'b0100111010010011100101001101010100110111;
	#t	xin=40'b0100110101010011011101001101110100111001;
	#t	xin=40'b0100111010010011010101001111010100110111;
	#t	xin=40'b0100111001010011000001001100110100110000;
	#t	xin=40'b0100110100010011011001001101110100110111;
	#t	xin=40'b0100110100010011011101001110100100110100;
	#t	xin=40'b0100111001010011101001001101100100110100;
	#t	xin=40'b0100110010010011000101001110110100111000;
	#t	xin=40'b0100110011010011101101001110000100111001;
	#t	xin=40'b0100110011010011100001001110100100111010;
	#t	xin=40'b0100110011010010110101001101110100111000;
	#t	xin=40'b0100110100010011000101001101100100110101;
	#t	xin=40'b0100111001010011001101001011110100110100;
	#t	xin=40'b0100111000010011011001001101010100110011;
	#t	xin=40'b0100110101010011100001001100100100110001;
	#t	xin=40'b0100110111010011011001001110100100110110;
	#t	xin=40'b0100111110010011011101001100110100110011;
	#t	xin=40'b0100110101010011010001001101000100110010;
	#t	xin=40'b0100110101010010111101001100010100101110;
	#t	xin=40'b0100110011010011010101001100110100110000;
	#t	xin=40'b0100110010010011000001001100100100101110;
	#t	xin=40'b0100110000010011001101001110010100110100;
	#t	xin=40'b0100101100010011000101001011010100110011;
	#t	xin=40'b0100110011010011010101001011010100110101;
	#t	xin=40'b0100110010010011001101001101010100110100;
	#t	xin=40'b0100110010010011001101001100110100111010;
	#t	xin=40'b0100110100010011011001001100010100110101;
	#t	xin=40'b0100110011010010111001001011110100101111;
	#t	xin=40'b0100110100010011001001001100100100110100;
	#t	xin=40'b0100110010010011001101001100100100101110;
	#t	xin=40'b0100110010010011001101001101010100111010;
	#t	xin=40'b0100110010010011001001001011010100110110;
	#t	xin=40'b0100110000010011011101001011100100101001;
	#t	xin=40'b0100101110010011000001001010010100101100;
	#t	xin=40'b0100110010010010111001001010110100101100;
	#t	xin=40'b0100111111010011101101001100010100101111;
	#t	xin=40'b0101010000010100011101001111110100110100;
	#t	xin=40'b0101010101010101010001010100110101010100;
	#t	xin=40'b0101100101010110101001011011100101110001;
	#t	xin=40'b0101111011011000010001100001010110001001;
	#t	xin=40'b0110001110011001010001100100110110010101;
	#t	xin=40'b0110010111011001110001100111010110011110;
	#t	xin=40'b0110011111011010010101101001000110100111;
	#t	xin=40'b0110100110011010011101101010000110101001;
	#t	xin=40'b0110101011011010111001101011100110101100;
	#t	xin=40'b0110110000011011000101101011100110110001;
	#t	xin=40'b0110110000011011000101101100010110110011;
	#t	xin=40'b0110110001011011001001101100110110110111;
	#t	xin=40'b0110110101011011010101101101100110110101;
	#t	xin=40'b0110110101011011011001101101110110111001;
	#t	xin=40'b0110110010011011001101101101100110110110;
	#t	xin=40'b0110101000011011000001101101000110110100;
	#t	xin=40'b0110100001011010100001101010010110101111;
	#t	xin=40'b0110001111011001011101100111100110011110;
	#t	xin=40'b0101110101010111111001100001110110000111;
	#t	xin=40'b0101010010010110000101011010100101101000;
	#t	xin=40'b0100110100010011101001001111110101000000;
	#t	xin=40'b0100100001010001110101000010110100001101;
	#t	xin=40'b0100001011001111110100111011110011011111;
	#t	xin=40'b0011111100001110001100110011110011010010;
	#t	xin=40'b0011011100001100111100110010110011010001;
	#t	xin=40'b0011010100001101011100110101010011010010;
	#t	xin=40'b0011011001001101100100110100100011010000;
	#t	xin=40'b0011011100001101110100110110100011010100;
	#t	xin=40'b0011011100001101101100111000010011011100;
	#t	xin=40'b0011011111001101110100111000110011011111;
	#t	xin=40'b0011100001001110001000111000000011100011;
	#t	xin=40'b0011100010001110011000111000110011011111;
	#t	xin=40'b0011100110001110010100111010100011101001;
	#t	xin=40'b0011100111001110011000111001100011101001;
	#t	xin=40'b0011110000001110111100111011110011101101;
	#t	xin=40'b0011110010001111000000111101110011110000;
	#t	xin=40'b0011101101001110011000111001110011110011;
	#t	xin=40'b0011101100001110110100111100010011110001;
	#t	xin=40'b0011101001001110110000111011000011110100;
	#t	xin=40'b0011110000001110101000111010110011101011;
	#t	xin=40'b0011110111001111010000111101010011110011;
	#t	xin=40'b0011110001001110111000111101000011110011;
	#t	xin=40'b0011101100001111011100111011010011110011;
	#t	xin=40'b0011101110001111000100111100010011110011;
	#t	xin=40'b0011101111001110110100111100000011110110;
	#t	xin=40'b0011101111001111101100111101000011110100;
	#t	xin=40'b0011110110001111101100111011100011101111;
	#t	xin=40'b0011111010001111001100111100100011110010;
	#t	xin=40'b0011110101001111001000111100010011101101;
	#t	xin=40'b0011110101001111001000111101010011110101;
	#t	xin=40'b0011101101001111000000111100110011111000;
	#t	xin=40'b0011101101001110111100111011000011101011;
	#t	xin=40'b0011110010001111000100111100010011101100;
	#t	xin=40'b0011110111001111000100111100010011110010;
	#t	xin=40'b0011110011001111000000111100110011101011;
	#t	xin=40'b0011110111001111001000111100110011110011;
	#t	xin=40'b0011110101001111011100111100000011110000;
	#t	xin=40'b0011110111001111011100111100100011110111;
	#t	xin=40'b0011111100001111101100111101100011111001;
	#t	xin=40'b0011110101001111000100111100100011110001;
	#t	xin=40'b0011110110001111000000111101100011110110;
	#t	xin=40'b0011110001001111010000111101010011110101;
	#t	xin=40'b0011110100001111100000111101010011110001;
	#t	xin=40'b0011111000001111110100111110100011110111;
	#t	xin=40'b0011111001001111100000111100010011110010;
	#t	xin=40'b0011110010001110111000111110010011110011;
	#t	xin=40'b0011110110001111010000111110000011110101;
	#t	xin=40'b0011111100001111111100111110000011111010;
	#t	xin=40'b0011111000001111110000111101100011110110;
	#t	xin=40'b0011111001001111011100111101110011110110;
	#t	xin=40'b0011110100010000000100111110000011110111;
	#t	xin=40'b0011111001001111101100111100110011110111;
	#t	xin=40'b0011111100001111101100111110010011110010;
	#t	xin=40'b0011110100001111100000111110000011110101;
	#t	xin=40'b0011111101001111100000111101110011111001;
	#t	xin=40'b0011111010001111011100111111100011111110;
	#t	xin=40'b0011111011001111100100111111100011111111;
	#t	xin=40'b0011111100001111111000111111000011111000;
	#t	xin=40'b0100000100001111011100111110110011111000;
	#t	xin=40'b0011111110001111101000111111000011110101;
	#t	xin=40'b0011111111001111110101000001000011111000;
	#t	xin=40'b0100000101010000000101000000010011111101;

	
    #t      $finish;
end
            
                            
endmodule                         
