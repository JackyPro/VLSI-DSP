//=======================================
// The Counter  (4-bit)
// IC Lab: Lab 03
// Date  : 2013.3.26
// vesion : v1.0
//=======================================

module counter(

clk,
rst,

dout

);


		
endmodule
    
    
    
    