//=======================================
// The Top module
// Design : yhchen
// Project: VLSI DSP Course
//=======================================


module Top(clk, rst, a0, a1, a2, a3, z0, z2, z4, z6);



endmodule

