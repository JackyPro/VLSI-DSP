module Top(en, up, clk, rst, dout);

input en, up;
input clk, rst;
output [15:0] dout;


endmodule