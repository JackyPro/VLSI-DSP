//=======================================
// The Top module
// Design : yhchen
// Project: VLSI DSP Course
//=======================================


module Top_1(clk, rst, a0, a1, a2, a3,a4,a5,a6,a7, z0,z1, z2,z3, z4,z5, z6,z7);

parameter w_i = 10;
parameter w_c = 12;
parameter w_o = w_i + w_c + 2;
parameter signed c1 = 12'b0111_1101_1000;//s7
parameter signed c2 = 12'b0111_0110_0100;//s6
parameter signed c3 = 12'b0110_1010_0111;
parameter signed c4 = 12'b0101_1010_1000;//s4
parameter signed c5 = 12'b0101_1100_1000;//s3
parameter signed c6 = 12'b0011_0000_1111;
parameter signed c7 = 12'b0001_1001_0000;//s1
/*
 c4=12'b0101_1010_1000
-s4=12'b1010_0101_1000
 s4=12'b0101_1010_1000
 c4=12'b0101_1010_1000

 c6=12'b0011_0000_1111
-s6=12'b1000_1001_1100
 s6=12'b0111_0110_0100
 c6=12'b0011_0000_1111

 c7=12'b0001_1001_0000
 s7=12'b0111_1101_1000
-s7=12'b1000_0010_1000
 c7=12'b0001_1001_0000

 c3=12'b0110_1010_0111
 s3=12'b0101_1100_1000
-s3=12'b1010_0011_1000
 c3=12'b0110_1010_0111

 c3=12'b0110_1010_0111
-s3=12'b1010_0011_1000
 s3=12'b0101_1100_1000
 c3=12'b0110_1010_0111

 c1=12'b0111_1101_1000
 s1=12'b0001_1001_0000
-s1=12'b1110_0111_0000
 c1=12'b0111_1101_1000
*/
input	signed [w_i-1:0]	a0, a2, a4, a6;
input	signed [w_i-1:0]	a1, a3, a5, a7;
input				clk, rst;
output	signed [w_o+1:0]	z0, z2, z4, z6;
output	signed [w_o+1:0]	z1, z3, z5, z7;
reg		signed [w_i-1:0]	aa0, aa2, aa4, aa6;
reg		signed [w_i-1:0]	aa1, aa3, aa5, aa7;
wire	signed [w_o-1:0]    zz00, zz01, zz02, zz03,
							zz40, zz41, zz42, zz43,
							zz20, zz21, zz22, zz23,
							zz60, zz61, zz62, zz63;
wire	signed [w_o-1:0]	zz10,zz11,zz30,zz31,zz50,zz51,zz70,zz71;
reg		signed [w_o+1:0]	z0, z2, z4, z6;
reg		signed [w_o+1:0]	z1, z3, z5, z7;

wire signed [w_i+1:0]	s0_01, s1_01, s2_01, s3_01,
						s0_76, s1_76, s2_76, s3_76,
						s0_32, s1_32, s2_32, s3_32,
						s0_45, s1_45, s2_45, s3_45,

						s0_30, s1_30, s2_30, s3_30,
						s0_47, s1_47, s2_47, s3_47,
						s0_12, s1_12, s2_12, s3_12,
						s0_65, s1_65, s2_65, s3_65,

						s0_03, s1_03, s2_03, s3_03,
						s0_74, s1_74, s2_74, s3_74,
						s0_21, s1_21, s2_21, s3_21,
						s0_56, s1_56, s2_56, s3_56;

//----- Input Reg ------//
always@(posedge clk) begin
	aa0 <= a0;
	aa2 <= a2;
	aa4 <= a4;
	aa6 <= a6;
	aa1 <= a1;
	aa3 <= a3;
	aa5 <= a5;
	aa7 <= a7;
end

//----- DA ------//
assign s0_01 = 0;
assign s1_01 = aa1;
assign s2_01 = aa0;
assign s3_01 = aa0 + aa1;

assign s0_76 = 0;
assign s1_76 = aa6;
assign s2_76 = aa7;
assign s3_76 = aa7 + aa6;

assign s0_32 = 0;
assign s1_32 = aa2;
assign s2_32 = aa3;
assign s3_32 = aa3 + aa2;

assign s0_45 = 0;
assign s1_45 = aa5;
assign s2_45 = aa4;
assign s3_45 = aa4 + aa5;

assign s0_30 = 0;
assign s1_30 = aa0;
assign s2_30 = aa3;
assign s3_30 = aa3 + aa0;

assign s0_47 = 0;
assign s1_47 = aa7;
assign s2_47 = aa4;
assign s3_47 = aa4 + aa7;

assign s0_12 = 0;
assign s1_12 = aa2;
assign s2_12 = aa1;
assign s3_12 = aa1 + aa2;

assign s0_65 = 0;
assign s1_65 = aa5;
assign s2_65 = aa6;
assign s3_65 = aa6 + aa5;

assign s0_03 = 0;
assign s1_03 = aa3;
assign s2_03 = aa0;
assign s3_03 = aa0 + aa3;

assign s0_74 = 0;
assign s1_74 = aa4;
assign s2_74 = aa7;
assign s3_74 = aa7 + aa4;

assign s0_21 = 0;
assign s1_21 = aa1;
assign s2_21 = aa2;
assign s3_21 = aa2 + aa1;

assign s0_56 = 0;
assign s1_56 = aa6;
assign s2_56 = aa5;
assign s3_56 = aa5 + aa6;

//----- Pipe -----//

//----- Add ------//
assign	zz40 = (s3_01<<3) + (s1_01<<4) + (s2_01<<5) + (s1_01<<6) + (s2_01<<7) + (s2_01<<8) + (s1_01<<9) + (s2_01<<10) + (s1_01<<11);
assign	zz41 = (s3_76<<3) + (s1_76<<4) + (s2_76<<5) + (s1_76<<6) + (s2_76<<7) + (s2_76<<8) + (s1_76<<9) + (s2_76<<10) + (s1_76<<11);
assign	zz42 = (s3_32<<3) + (s1_32<<4) + (s2_32<<5) + (s1_32<<6) + (s2_32<<7) + (s2_32<<8) + (s1_32<<9) + (s2_32<<10) + (s1_32<<11);
assign	zz43 = (s3_45<<3) + (s1_45<<4) + (s2_45<<5) + (s1_45<<6) + (s2_45<<7) + (s2_45<<8) + (s1_45<<9) + (s2_45<<10) + (s1_45<<11);

assign	zz00 = (s3_01<<3) + (s3_01<<5) + (s3_01<<7) + (s3_01<<8) + (s3_01<<10);
assign	zz01 = (s3_76<<3) + (s3_76<<5) + (s3_76<<7) + (s3_76<<8) + (s3_76<<10);
assign	zz02 = (s3_32<<3) + (s3_32<<5) + (s3_32<<7) + (s3_32<<8) + (s3_32<<10);
assign	zz03 = (s3_45<<3) + (s3_45<<5) + (s3_45<<7) + (s3_45<<8) + (s3_45<<10);

assign	zz60 =  s2_01 + (s2_01<<1) + (s3_01<<2) + (s3_01<<3) + (s1_01<<4) + (s1_01<<7) + (s2_01<<8) + (s2_01<<9) + (s1_01<<11);
assign	zz61 =  s2_76 + (s2_76<<1) + (s3_76<<2) + (s3_76<<3) + (s1_76<<4) + (s1_76<<7) + (s2_76<<8) + (s2_76<<9) + (s1_76<<11);
assign	zz62 =  s2_32 + (s2_32<<1) + (s3_32<<2) + (s3_32<<3) + (s1_32<<4) + (s1_32<<7) + (s2_32<<8) + (s2_32<<9) + (s1_32<<11);
assign	zz63 =  s2_45 + (s2_45<<1) + (s3_45<<2) + (s3_45<<3) + (s1_45<<4) + (s1_45<<7) + (s2_45<<8) + (s2_45<<9) + (s1_45<<11);

assign	zz20 =  s1_01 + (s1_01<<1) + (s3_01<<2) + (s1_01<<3) + (s2_01<<5) + (s2_01<<6) + (s3_01<<8) + (s3_01<<9) + (s2_01<<10);
assign	zz21 =  s1_76 + (s1_76<<1) + (s3_76<<2) + (s1_76<<3) + (s2_76<<5) + (s2_76<<6) + (s3_76<<8) + (s3_76<<9) + (s2_76<<10);
assign	zz22 =  s1_32 + (s1_32<<1) + (s3_32<<2) + (s1_32<<3) + (s2_32<<5) + (s2_32<<6) + (s3_32<<8) + (s3_32<<9) + (s2_32<<10);
assign	zz23 =  s1_45 + (s1_45<<1) + (s3_45<<2) + (s1_45<<3) + (s2_45<<5) + (s2_45<<6) + (s3_45<<8) + (s3_45<<9) + (s2_45<<10);


assign  zz10 =  (s1_30<<3) + (s3_30<<4) + (s1_30<<6) + (s3_30<<7) + (s3_30<<8) + (s1_30<<9) + (s1_30<10)
             + s2_12 + (s2_12<<1) + (s2_12<<2) + (s1_12<<3) + (s2_12<<5) + (s1_12<<6) + (s3_12<<7) + (s1_12<<8) + (s2_12<<9) + (s3_12<<10);
assign  zz11 =  (s1_47<<3) + (s3_47<<4) + (s1_47<<6) + (s3_47<<7) + (s3_47<<8) + (s1_47<<9) + (s1_47<10)
             + s2_65 + (s2_65<<1) + (s2_65<<2) + (s1_65<<3) + (s2_65<<5) + (s1_65<<6) + (s3_65<<7) + (s1_65<<8) + (s2_65<<9) + (s3_65<<10);

assign  zz70 =  (s2_30<<3) + (s1_30<<4) + (s2_30<<5) + (s1_30<<7) + (s1_30<<8) + (s2_30<<11) 
             + s1_12 + (s1_12<<1) + (s1_12<<2) + (s2_12<<3) + (s2_12<<4) + (s3_12<<5) + (s1_12<<7) + (s3_12<<9) + (s1_12<<10) + (s2_12<<11); 
assign  zz71 =  (s2_47<<3) + (s1_47<<4) + (s2_47<<5) + (s1_47<<7) + (s1_47<<8) + (s2_47<<11) 
             + s1_65 + (s1_65<<1) + (s1_65<<2) + (s2_65<<3) + (s2_65<<4) + (s3_65<<5) + (s1_65<<7) + (s3_65<<9) + (s1_65<<10) + (s2_65<<11); 

assign  zz30 =  s2_03 + (s2_03<<1) + (s2_03<<2) + (s1_03<<3) + (s1_03<<4) + (s3_03<<5) + (s2_03<<7) + (s3_03<<9) + (s2_03<<10) + (s1_03<<11)
             -( (s2_21<<3) + (s3_21<<4) + (s2_21<<6) + (s3_21<<7) + (s3_21<<8) + (s2_21<<9) + (s2_21<<10) );
assign  zz31 =  s2_74 + (s2_74<<1) + (s2_74<<2) + (s1_74<<3) + (s1_74<<4) + (s3_74<<5) + (s2_74<<7) + (s3_74<<9) + (s2_74<<10) + (s1_74<<11)
             -( (s2_56<<3) + (s3_56<<4) + (s2_56<<6) + (s3_56<<7) + (s3_56<<8) + (s2_56<<9) + (s2_56<<10) );

assign  zz50 =  s1_03 + (s1_03<<1) + (s1_03<<2) + (s2_03<<3) + (s1_03<<5) + (s2_03<<6) + (s3_03<<7) + (s2_03<<8) + (s1_03<<9) + (s3_03<<10)
             -( (s1_21<<3) + (s3_21<<4) + (s2_21<<5) + (s3_21<<6) + (s1_21<<7) + (s1_21<<8) +(s3_21<<9) + (s3_21<<10) + (s2_21<<11) );
assign  zz51 =  s1_74 + (s1_74<<1) + (s1_74<<2) + (s2_74<<3) + (s1_74<<5) + (s2_74<<6) + (s3_74<<7) + (s2_74<<8) + (s1_74<<9) + (s3_74<<10)
             -( (s1_56<<3) + (s3_56<<4) + (s2_56<<5) + (s3_56<<6) + (s1_56<<7) + (s1_56<<8) +(s3_56<<9) + (s3_56<<10) + (s2_56<<11) );


//----- Output Reg ------//
always@(posedge clk) begin
	z0 <= zz00+zz01+zz02+zz03;
    z1 <= zz10-zz11;
	z2 <= zz20+zz21-zz22-zz23;
    z3 <= zz30-zz31;
	z4 <= zz40+zz41+zz42+zz43;
    z5 <= zz50-zz51;
	z6 <= zz60+zz61-zz62-zz63;
    z7 <= zz70-zz71;
end

endmodule

